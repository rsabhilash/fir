module carry_select_adder #(
parameter IN_DATAWIDTH = 8 ,
parameter OUT_DATAWIDTH = IN_DATAWIDTH+1
)
(
input [IN_DATAWIDTH-1:0] in1 ,
input [IN_DATAWIDTH-1:0] in2 ,
output [OUT_DATAWIDTH-1:0] out
);

endmodule


